

package chm_tb_cor_pkg;

    import uvm_pkg::*;
    import uvme_cv32e20_pkg::*;
    import uvmt_cv32e20_pkg::*;

    `include "uvm_macros.svh"

    `include "chm_tb_cor_test.sv"

endpackage
